----------------------------------------------------------------------------------
-- COPYRIGHT 2019 Jes�s Eduardo M�ndez Rosales
--This program is free software: you can redistribute it and/or modify
--it under the terms of the GNU General Public License as published by
--the Free Software Foundation, either version 3 of the License, or
--(at your option) any later version.
--
--This program is distributed in the hope that it will be useful,
--but WITHOUT ANY WARRANTY; without even the implied warranty of
--MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--GNU General Public License for more details.
--
--You should have received a copy of the GNU General Public License
--along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--
--							LIBRER�A LCD
--
-- Descripci�n: Con �sta librer�a podr�s implementar c�digos para una LCD 16x2 de manera
-- f�cil y r�pida, con todas las ventajas de utilizar una FPGA.
--
-- Caracter�sticas:
-- 
--	Los comandos que puedes utilizar son los siguientes:
--
-- LCD_INI() -> Inicializa la lcd.
--		 			 NOTA: Dentro de los par�ntesis poner un vector de 2 bits para encender o apagar
--					 		 el cursor y activar o desactivar el parpadeo.
--
--		"1x" -- Cursor ON
--		"0x" -- Cursor OFF
--		"x1" -- Parpadeo ON
--		"x0" -- Parpadeo OFF
--
--   Por ejemplo: LCD_INI("10") -- Inicializar LCD con cursor encendido y sin parpadeo 
--	
--			
-- CHAR() -> Manda una letra may�scula o min�scula
--
--				 IMPORTANTE: 1) Debido a que VHDL no es sensible a may�sculas y min�sculas, si se quiere
--								    escribir una letra may�scula se debe escribir una "M" antes de la letra.
--								 2) Si se quiere escribir la letra "S" may�scula, se declara "MAS"
--											
-- 	Por ejemplo: CHAR(A)  -- Escribe en la LCD la letra "a"
--						 CHAR(MA) -- Escribe en la LCD la letra "A"	
--						 CHAR(S)	 -- Escribe en la LCD la letra "s"
--						 CHAR(MAS)	 -- Escribe en la LCD la letra "S"	
--	
--
-- POS() -> Escribir en la posici�n que se indique.
--				NOTA: Dentro de los par�ntesis se dene poner la posici�n de la LCD a la que se quiere ir, empezando
--						por el rengl�n seguido de la posici�n vertical, ambos n�meros separados por una coma.
--		
--		Por ejemplo: POS(1,2) -- Manda cursor al rengl�n 1, poscici�n 2
--						 POS(2,4) -- Manda cursor al rengl�n 2, poscici�n 4		
--
--
-- CHAR_ASCII() -> Escribe un caracter a partir de su c�digo en ASCII
--						 NOTA: Dentro de los parentesis escribir x"(n�mero hex.)"
--
--		Por ejemplo: CHAR_ASCII(x"40") -- Escribe en la LCD el caracter "@"
--
--
-- CODIGO_FIN() -> Finaliza el c�digo. 
--						 NOTA: Dentro de los par�ntesis poner cualquier n�mero: 1,2,3,4...,8,9.
--
--
-- BUCLE_INI() -> Indica el inicio de un bucle. 
--						NOTA: Dentro de los par�ntesis poner cualquier n�mero: 1,2,3,4...,8,9.
--
--
-- BUCLE_FIN() -> Indica el final del bucle.
--						NOTA: Dentro de los par�ntesis poner cualquier n�mero: 1,2,3,4...,8,9.
--
--
-- INT_NUM() -> Escribe en la LCD un n�mero entero.
--					 NOTA: Dentro de los par�ntesis poner s�lo un n�mero que vaya del 0 al 9,
--						    si se quiere escribir otro n�mero entero se tiene que volver
--							 a llamar la funci�n
--
--
-- CREAR_CHAR() -> Funci�n que crea el caracter dise�ado previamente en "CARACTERES_ESPECIALES.vhd"
--                 NOTA: Dentro de los par�ntesis poner el nombre del caracter dibujado (CHAR1,CHAR2,CHAR3,..,CHAR8)
--								 
--
-- CHAR_CREADO() -> Escribe en la LCD el caracter creado por medio de la funci�n "CREAR_CHAR()"
--						  NOTA: Dentro de los par�ntesis poner el nombre del caracter creado.
--
--     Por ejemplo: 
--
--				Dentro de CARACTERES_ESPECIALES.vhd se dibujan los caracteres personalizados utilizando los vectores 
--				"CHAR_1", "CHAR_2","CHAR_3",...,"CHAR_7","CHAR_8"
--
--								 '1' => [#] - Se activa el pixel de la matr�z.
--                       '0' => [ ] - Se desactiva el pixel de la matriz.
--
-- 			Si se quiere crear el				Entonces CHAR_1 queda de la siguiente
--				siguiente caracter:					manera:
--												
--				  1  2  3  4  5						CHAR_1 <=
--  		  1 [ ][ ][ ][ ][ ]							"00000"&			
-- 		  2 [ ][ ][ ][ ][ ]							"00000"&			  
-- 		  3 [ ][#][ ][#][ ]							"01010"&   		  
-- 		  4 [ ][ ][ ][ ][ ]		=====>			"00000"&			   
-- 		  5 [#][ ][ ][ ][#]							"10001"&          
-- 		  6 [ ][#][#][#][ ]							"01110"&			  
-- 		  7 [ ][ ][ ][ ][ ]							"00000"&			  
-- 		  8 [ ][ ][ ][ ][ ]							"00000";			
--
--		
--			Como el caracter se cre� en el vector "CHAR_1",entonces se escribe en las funci�nes como "CHAR1"
--			
--			CREAR_CHAR(CHAR1)  -- Crea el caracter personalizado (CHAR1)
--			CHAR_CREADO(CHAR1) -- Muestra en la LCD el caracter creado (CHAR1)		
--
-- 
--
-- LIMPIAR_PANTALLA() -> Manda a limpiar la LCD.
--								 NOTA: �sta funci�n se activa poniendo dentro de los par�ntesis
--										 un '1' y se desactiva con un '0'. 
--
--		Por ejemplo: LIMPIAR_PANTALLA('1') -- Limpiar pantalla est� activado.
--						 LIMPIAR_PANTALLA('0') -- Limpiar pantalla est� desactivado.
--
--
--	Con los puertos de entrada "CORD" y "CORI" se hacen corrimientos a la derecha y a la
--	izquierda respectivamente. NOTA: La velocidad del corrimiento se puede cambiar 
-- modificando la variable "DELAY_COR".
--
-- Algunas funci�nes generan un vector ("BLCD") cuando se termin� de ejecutar dicha funci�n y
--	que puede ser utilizado como una bandera, el vector solo dura un ciclo de instruccion.
--	   
--		LCD_INI() ---------- BLCD <= x"01"
--		CHAR() ------------- BLCD <= x"02"
--		POS() -------------- BLCD <= x"03"
-- 	INT_NUM() ---------- BLCD <= x"04"
--	   CHAR_ASCII() ------- BLCD <= x"05"
--	   BUCLE_INI() -------- BLCD <= x"06"
--		BUCLE_FIN() -------- BLCD <= x"07"
--		LIMPIAR_PANTALLA() - BLCD <= x"08"
--	   CREAR_CHAR() ------- BLCD <= x"09"
--	 	CHAR_CREADO() ------ BLCD <= x"0A"
--
--
--		�IMPORTANTE!
--		
--		1) Se deber� especificar el n�mero de instrucciones en la constante "NUM_INSTRUCCIONES". El valor 
--			de la �ltima instrucci�n es el que se colocar�
--		2) En caso de utilizar a la librer�a como TOP del dise�o, se deber� comentar el puerto gen�rico y 
--			descomentar la constante "FPGA_CLK" para especificar la frecuencia de reloj.
--		3) Cada funci�n se acompa�a con " INST(NUM) <= <FUNCI�N> " como lo muestra en el c�digo
-- 		demostrativo.
--
--
--                C�DIGO DEMOSTRATIVO
--
--		CONSTANT NUM_INSTRUCCIONES : INTEGER := 7;
--
-- 	INST(0) <= LCD_INI("11"); 		-- INICIALIZAMOS LCD, CURSOR A HOME, CURSOR ON, PARPADEO ON.
-- 	INST(1) <= POS(1,1);				-- EMPEZAMOS A ESCRIBIR EN LA LINEA 1, POSICI�N 1
-- 	INST(2) <= CHAR(MH);				-- ESCRIBIMOS EN LA LCD LA LETRA "h" MAYUSCULA
-- 	INST(3) <= CHAR(O);			
-- 	INST(4) <= CHAR(L);
-- 	INST(5) <= CHAR(A);
-- 	INST(6) <= CHAR_ASCII(x"21"); -- ESCRIBIMOS EL CARACTER "!"
-- 	INST(7) <= CODIGO_FIN(1);	   -- FINALIZAMOS EL CODIGO
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE WORK.COMANDOS_LCD_REVD.ALL;

entity LIB_LCD_INTESC_REVD is

GENERIC(
			FPGA_CLK : INTEGER := 50_000_000
);


PORT(CLK: IN STD_LOGIC;

-----------------------------------------------------
------------------PUERTOS DE LA LCD------------------
	  RS 		  : OUT STD_LOGIC;							--
	  RW		  : OUT STD_LOGIC;							--
	  ENA 	  : OUT STD_LOGIC;							--
	  DATA_LCD : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);  --
-----------------------------------------------------
-----------------------------------------------------
	  
	  
-----------------------------------------------------------
--------------ABAJO ESCRIBE TUS PUERTOS--------------------	
	 	gripper: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		base : IN STD_LOGIC_VECTOR(6 DOWNTO 0)
-----------------------------------------------------------
-----------------------------------------------------------

	  );

end LIB_LCD_INTESC_REVD;

architecture Behavioral of LIB_LCD_INTESC_REVD is


CONSTANT NUM_INSTRUCCIONES : INTEGER := 36; 	--INDICAR EL N�MERO DE INSTRUCCIONES PARA LA LCD


--------------------------------------------------------------------------------
-------------------------SE�ALES DE LA LCD (NO BORRAR)--------------------------
																										--
component PROCESADOR_LCD_REVD is																--
																										--
GENERIC(																								--
			FPGA_CLK : INTEGER := 50_000_000;												--
			NUM_INST : INTEGER := 1																--
);																										--
																										--
PORT( CLK 				 : IN  STD_LOGIC;														--
	   VECTOR_MEM 		 : IN  STD_LOGIC_VECTOR(8  DOWNTO 0);							--
	   C1A,C2A,C3A,C4A : IN  STD_LOGIC_VECTOR(39 DOWNTO 0);							--
	   C5A,C6A,C7A,C8A : IN  STD_LOGIC_VECTOR(39 DOWNTO 0);							--
	   RS 				 : OUT STD_LOGIC;														--
	   RW 				 : OUT STD_LOGIC;														--
	   ENA 				 : OUT STD_LOGIC;														--
	   BD_LCD 			 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);			         	--
	   DATA 				 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);							--
	   DIR_MEM 			 : OUT INTEGER RANGE 0 TO NUM_INSTRUCCIONES					--
	);																									--
																										--
end component PROCESADOR_LCD_REVD;															--
																										--
COMPONENT CARACTERES_ESPECIALES_REVD is													--
																										--
PORT( C1,C2,C3,C4 : OUT STD_LOGIC_VECTOR(39 DOWNTO 0);								--
		C5,C6,C7,C8 : OUT STD_LOGIC_VECTOR(39 DOWNTO 0)									--
	 );																								--
																										--
end COMPONENT CARACTERES_ESPECIALES_REVD;													--
																										--
CONSTANT CHAR1 : INTEGER := 1;																--
CONSTANT CHAR2 : INTEGER := 2;																--
CONSTANT CHAR3 : INTEGER := 3;																--
CONSTANT CHAR4 : INTEGER := 4;																--
CONSTANT CHAR5 : INTEGER := 5;																--
CONSTANT CHAR6 : INTEGER := 6;																--
CONSTANT CHAR7 : INTEGER := 7;																--
CONSTANT CHAR8 : INTEGER := 8;																--
																										--
type ram is array (0 to  NUM_INSTRUCCIONES) of std_logic_vector(8 downto 0); 	--
signal INST : ram := (others => (others => '0'));										--
																										--
signal blcd 			  : std_logic_vector(7 downto 0):= (others => '0');		--																										
signal vector_mem 	  : STD_LOGIC_VECTOR(8  DOWNTO 0) := (others => '0');		--
signal c1s,c2s,c3s,c4s : std_logic_vector(39 downto 0) := (others => '0');		--
signal c5s,c6s,c7s,c8s : std_logic_vector(39 downto 0) := (others => '0'); 	--
signal dir_mem 		  : integer range 0 to NUM_INSTRUCCIONES := 0;				--
																										--
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
---------------------------AGREGA TUS SE�ALES AQU�------------------------------
CONSTANT ABRIENDO : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
CONSTANT CERRANDO : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
CONSTANT GIRODER : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
CONSTANT GIROIZQ : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
CONSTANT DETENIDO : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
SIGNAL ESTADO_GRIPPER : STD_LOGIC_VECTOR (1 DOWNTO 0);
SIGNAL ESTADO_BASE : STD_LOGIC_VECTOR (1 DOWNTO 0);
SIGNAL P_GRIPPER : STD_LOGIC_VECTOR(63 downto 0);
SIGNAL P_BASE : STD_LOGIC_VECTOR(63 downto 0);
SIGNAL CONT_GB : INTEGER;
SIGNAL SAMPLED_GRIPPER : STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL SAMPLED_BASE : STD_LOGIC_VECTOR(6 DOWNTO 0);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------


begin


---------------------------------------------------------------
-------------------COMPONENTES PARA LCD------------------------
																				 --
u1: PROCESADOR_LCD_REVD													 --
GENERIC map( FPGA_CLK => FPGA_CLK,									 --
				 NUM_INST => NUM_INSTRUCCIONES )						 --
																				 --
PORT map( CLK,VECTOR_MEM,C1S,C2S,C3S,C4S,C5S,C6S,C7S,C8S,RS, --
			 RW,ENA,BLCD,DATA_LCD, DIR_MEM );						 --
																				 --
U2 : CARACTERES_ESPECIALES_REVD 										 --
PORT MAP( C1S,C2S,C3S,C4S,C5S,C6S,C7S,C8S );				 		 --
																				 --
VECTOR_MEM <= INST(DIR_MEM);											 --
																				 --
---------------------------------------------------------------
---------------------------------------------------------------


-------------------------------------------------------------------
---------------ESCRIBE TU C�DIGO PARA LA LCD-----------------------

 	INST(0) <= LCD_INI("00"); 		-- INICIALIZAMOS LCD, CURSOR A HOME, CURSOR ON, PARPADEO ON.
 	INST(1) <= POS(1,1);				-- EMPEZAMOS A ESCRIBIR EN LA LINEA 1, POSICI�N 1
	
	-- 1234567890123456	1234567890123456	1234567890123456
	-- Gripper:ABRIENDO	Gripper:CERRANDO	Gripper:DETENIDO
	-- Base:***GIRO*DER	Base:***GIRO*IZQ	Base:***DETENIDO
	
	INST(2) <= CHAR(MG);				--G
	INST(3) <= CHAR(R);				--r
	INST(4) <= CHAR(I);				--i
	INST(5) <= CHAR(P);				--p
	INST(6) <= CHAR(P);				--p
	INST(7) <= CHAR(E);				--e
	INST(8) <= CHAR(R);				--r
	INST(9) <= CHAR_ASCII(x"3A"); --:
	INST(10) <= POS(2,1);
	INST(11) <= CHAR(MB);			--B
	INST(12) <= CHAR(a);				--a
	INST(13) <= CHAR(s);				--s
	INST(14) <= CHAR(e);				--e
	INST(15) <= CHAR_ASCII(x"3A");--:
	
	INST(16) <= BUCLE_INI(1);
	INST(17) <= POS(1,9);

	INST(18) <= CHAR_ASCII(P_GRIPPER(63 downto 56));	--A C D
	INST(19) <= CHAR_ASCII(P_GRIPPER(55 downto 48));	--B E E
	INST(20) <= CHAR_ASCII(P_GRIPPER(47 downto 40));	--R R T
	INST(21) <= CHAR_ASCII(P_GRIPPER(39 downto 32));	--I R E
	INST(22) <= CHAR_ASCII(P_GRIPPER(31 downto 24));	--E A N
	INST(23) <= CHAR_ASCII(P_GRIPPER(23 downto 16));	--N N I
	INST(24) <= CHAR_ASCII(P_GRIPPER(15 downto 8));		--D D D
	INST(25) <= CHAR_ASCII(P_GRIPPER(7 downto 0));		--O O O

	INST(26) <= POS(2,9);

	INST(27) <= CHAR_ASCII(P_BASE(63 downto 56));	--G G D
	INST(28) <= CHAR_ASCII(P_BASE(55 downto 48));	--I I E
	INST(29) <= CHAR_ASCII(P_BASE(47 downto 40));	--R R T
	INST(30) <= CHAR_ASCII(P_BASE(39 downto 32));	--O O E
	INST(31) <= CHAR_ASCII(P_BASE(31 downto 24));	--    N
	INST(32) <= CHAR_ASCII(P_BASE(23 downto 16));	--D I I
	INST(33) <= CHAR_ASCII(P_BASE(15 downto 8));		--E Z D
	INST(34) <= CHAR_ASCII(P_BASE(7 downto 0));		--R Q O
	
	INST(35) <= BUCLE_FIN(1);
	
 	INST(36) <= CODIGO_FIN(1);	   -- FINALIZAMOS EL CODIGO

-------------------------------------------------------------------
-------------------------------------------------------------------




-------------------------------------------------------------------
--------------------ESCRIBE TU C�DIGO DE VHDL----------------------
PROCESS(ESTADO_GRIPPER) BEGIN
		CASE ESTADO_GRIPPER IS
		WHEN ABRIENDO => P_GRIPPER <= (X"41"&X"42"&X"52"&X"49"&X"45"&X"4e"&X"44"&X"4f"); -- ABRIENDO
		WHEN CERRANDO => P_GRIPPER <= (X"43"&X"45"&X"52"&X"52"&X"41"&X"4e"&X"44"&X"4f"); -- CERRANDO
		WHEN OTHERS => P_GRIPPER <= (X"44"&X"45"&X"54"&X"45"&X"4e"&X"49"&X"44"&X"4f"); -- DETENIDO
		END CASE;
END PROCESS;

PROCESS(ESTADO_BASE) BEGIN
	CASE ESTADO_BASE IS
		WHEN GIRODER => P_BASE <= (X"47"&X"49"&X"52"&X"4f"&X"20"&X"44"&X"45"&X"52"); -- GIRO DER
		WHEN GIROIZQ => P_BASE <= (X"47"&X"49"&X"52"&X"4f"&X"20"&X"49"&X"5a"&X"51"); -- CERRANDO
		WHEN OTHERS => P_BASE <= (X"44"&X"45"&X"54"&X"45"&X"4e"&X"49"&X"44"&X"4f"); -- DETENIDO
		END CASE;
END PROCESS;

PROCESS(CLK, GRIPPER, BASE) BEGIN
	IF( CLK'EVENT AND CLK='1' ) THEN
		IF( CONT_GB = 24_999_999 ) THEN 
			CONT_GB <= 0;
			IF( GRIPPER < SAMPLED_GRIPPER ) THEN ESTADO_GRIPPER <= CERRANDO;
			ELSIF( GRIPPER > SAMPLED_GRIPPER ) THEN ESTADO_GRIPPER <= ABRIENDO;
			ELSE ESTADO_GRIPPER <= DETENIDO;
			END IF;
			IF( BASE > SAMPLED_BASE ) THEN ESTADO_BASE <= GIROIZQ;
			ELSIF( BASE < SAMPLED_BASE ) THEN ESTADO_BASE <= GIRODER;
			ELSE ESTADO_BASE <= DETENIDO;
			END IF;
		ELSE
			CONT_GB <= CONT_GB + 1;
			IF(CONT_GB = 0) THEN 
				SAMPLED_GRIPPER <= GRIPPER;
				SAMPLED_BASE <= BASE;
			END IF;
		END IF;
	END IF;
END PROCESS;

-------------------------------------------------------------------
-------------------------------------------------------------------





end Behavioral;

