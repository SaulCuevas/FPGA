-- INSTITUTO POLITECNICO NACIONAL
-- 				UPIITA
-- AUTORES: SAUL CUEVAS MORALES
-- 			ALEXIS GONZALEZ ZUNIGA
-- SENSORES E INICIO
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BOTON is
port(
		CLK : IN STD_LOGIC; 							--RELOJ DE 50MHz
		ENABLE : IN STD_LOGIC; 						--BOTON DE ENCENDIDO / APAGADO 
		
		SENSD : IN STD_LOGIC;						--SENSOR DE LA DERECHA
		SENSI : IN STD_LOGIC;						--SENSOR DE LA IZQUIERDA
		
		SENTIDO : INOUT STD_LOGIC						--BIT DETERMINANTE DEL SENTIDO "1" -> DERECHA, "0" -> IZQUIERDA
);	
end BOTON;

architecture Behavioral of BOTON is

begin	
	PROCESS(CLK, ENABLE, SENSD, SENSI) BEGIN
		IF(CLK'event AND CLK = '1' AND ENABLE = '1') THEN
			IF(SENSD = '1') THEN SENTIDO <= '0';
			ELSIF (SENSI = '1') THEN SENTIDO <= '1';
			ELSIF (SENTIDO /= '1' AND SENTIDO /= '0') THEN SENTIDO <= '1';
			ELSE SENTIDO <= SENTIDO;
			END IF;
		END IF;
	END PROCESS;
end Behavioral;

