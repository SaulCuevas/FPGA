----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SEMAFOROS is
    Port ( CLK			  : in	STD_LOGIC; 		--50MHz
			  SEMAFORO_NS : out  STD_LOGIC_VECTOR(2 DOWNTO 0);
           SEMAFORO_EO : out  STD_LOGIC_VECTOR(2 DOWNTO 0);
           FOTORESISTENCIA : in  STD_LOGIC;
           PEATONAL_COLS :	out	STD_LOGIC_VECTOR(7 DOWNTO 0); 	--COLUMNAS DE LA MATRIZ DE LEDS
			  PEATONAL_FILS :	inout  	STD_LOGIC_VECTOR(15 DOWNTO 0); 	--FILAS DE LA MATRIZ DE LEDS
			  BOCINA : 			out 	STD_LOGIC);	--PARA MENSAJES DE VOZ
           --RELOJ_1HZ : in  STD_LOGIC);			--RELOJ EXTERNO
end SEMAFOROS;

architecture Behavioral of SEMAFOROS is
SIGNAL RELOJ_1HZ : STD_LOGIC;
SIGNAL RELOJ_80HZ : STD_LOGIC;
SIGNAL RELOJ_240HZ : STD_LOGIC;
SIGNAL RELOJ_960HZ : STD_LOGIC;

SIGNAL FILAS : INTEGER RANGE 1 TO 16:=1;
SIGNAL ANIMACION : STD_LOGIC_VECTOR(1 DOWNTO 0);

signal conta : integer range 1 to 25_000_000:=1; 
signal conta_ulti : integer :=25_000_000;

signal conta_1 : integer range 1 to 26_042:=1; 
signal conta_ulti_1 : integer :=26_042;

signal conta_2 : integer range 1 to 312_500:=1; 
signal conta_ulti_2 : integer :=312_500;

signal conta_3 : integer range 1 to 104_167:=1; 
signal conta_ulti_3 : integer :=104_167;

SIGNAL CONTADOR : INTEGER RANGE 0 TO 29:=0;
SIGNAL MS_500 : INTEGER RANGE 1 TO 12_500_000:=1;
begin

	--GENERANDO LA SENAL DE 1HZ----------
	process (CLK) begin
		if rising_edge(CLK) then
			if (conta = conta_ulti) then
				RELOJ_1HZ <= NOT(RELOJ_1HZ);
				conta <= 1;
			else
				conta <= conta + 1;
			end if;
		end if;
	end process;
	
	--GENERANDO LA SENAL DE 960HZ----------
	process (CLK) begin
		if rising_edge(CLK) then
			if (conta_1 = conta_ulti_1) then
				RELOJ_960HZ <= NOT(RELOJ_960HZ);
				conta_1 <= 1;
			else
				conta_1 <= conta_1 + 1;
			end if;
		end if;
	end process;

	--GENERANDO LA SENAL DE 80HZ----------
	process (CLK) begin
		if rising_edge(CLK) then
			if (conta_2 = conta_ulti_2) then
				RELOJ_80HZ <= NOT(RELOJ_80HZ);
				conta_2 <= 1;
			else
				conta_2 <= conta_2 + 1;
			end if;
		end if;
	end process;

	--GENERANDO LA SENAL DE 240HZ----------
	process (CLK) begin
		if rising_edge(CLK) then
			if (conta_3 = conta_ulti_3) then
				RELOJ_240HZ <= NOT(RELOJ_240HZ);
				conta_3 <= 1;
			else
				conta_3 <= conta_3 + 1;
			end if;
		end if;
	end process;
	
	--PROCESO PARA EL CONTADOR--------------------
	PROCESS(CLK, RELOJ_1HZ, CONTADOR) BEGIN
		IF RISING_EDGE(CLK) THEN
			IF CONTADOR <= 5 AND CONTADOR >= 11 THEN
				IF MS_500 = 12_500_000 THEN 
					CONTADOR <= CONTADOR + 1;
					MS_500 <= 1;
				ELSE MS_500 <= MS_500 + 1;
				END IF;
			ELSIF CONTADOR <= 20 AND CONTADOR >= 26 THEN
				IF MS_500 = 12_500_000 THEN 
					CONTADOR <= CONTADOR + 1;
					MS_500 <= 1;
				ELSE MS_500 <= MS_500 + 1;
				END IF;
			ELSE 
				IF RISING_EDGE(RELOJ_1HZ) THEN
					CONTADOR <= CONTADOR + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	--ANIMACION DE MATRIZ DE LEDS-----------
	PROCESS(CLK, CONTADOR) BEGIN
		IF RISING_EDGE(CLK) THEN
			IF CONTADOR >= 15 THEN ANIMACION <= "00";
			ELSIF CONTADOR >= 0 AND CONTADOR < 12 THEN 
				IF RISING_EDGE(RELOJ_80HZ) THEN
					ANIMACION <= ANIMACION + 1;
				END IF;
			ELSIF CONTADOR >= 12 AND CONTADOR < 15 THEN
				IF RISING_EDGE(RELOJ_240HZ) THEN
					ANIMACION <= ANIMACION + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	--SEMAFOROS-----------------------------
	PROCESS(CLK, FOTORESISTENCIA, CONTADOR) BEGIN
		IF RISING_EDGE(CLK) THEN
			IF FOTORESISTENCIA = '0' THEN --MODO NORMAL
				CASE CONTADOR IS
					WHEN 0 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 1 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 2 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 3 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 4 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 5 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 6 => SEMAFORO_NS <= "000"; SEMAFORO_EO <= "001";
					WHEN 7 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 8 => SEMAFORO_NS <= "000"; SEMAFORO_EO <= "001";
					WHEN 9 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 10 => SEMAFORO_NS <= "000"; SEMAFORO_EO <= "001";
					WHEN 11 => SEMAFORO_NS <= "100"; SEMAFORO_EO <= "001";
					WHEN 12 => SEMAFORO_NS <= "010"; SEMAFORO_EO <= "001";
					WHEN 13 => SEMAFORO_NS <= "010"; SEMAFORO_EO <= "001";
					WHEN 14 => SEMAFORO_NS <= "010"; SEMAFORO_EO <= "001";
					WHEN 15 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 16 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 17 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 18 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 19 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 20 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 21 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "000";
					WHEN 22 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 23 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "000";
					WHEN 24 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 25 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "000";
					WHEN 26 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "100";
					WHEN 27 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "010";
					WHEN 28 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "010";
					WHEN 29 => SEMAFORO_NS <= "001"; SEMAFORO_EO <= "010";
					WHEN OTHERS => SEMAFORO_NS <= "000"; SEMAFORO_EO <= "000";
				END CASE;
			ELSE --MODO NORMAL
			END IF;
		END IF;
	END PROCESS;
	
	--CAMBIO DE FILA----------------------------------------------
	PROCESS(CLK, RELOJ_960HZ, FILAS) BEGIN
		IF RISING_EDGE(CLK) THEN
			IF RISING_EDGE(RELOJ_960HZ) THEN
				FILAS <= FILAS + 1;
				CASE FILAS IS
					WHEN 1	 => PEATONAL_FILS <= NOT("0000000000000001");
					WHEN 2	 => PEATONAL_FILS <= NOT("0000000000000010");
					WHEN 3	 => PEATONAL_FILS <= NOT("0000000000000100");
					WHEN 4	 => PEATONAL_FILS <= NOT("0000000000001000");
					WHEN 5	 => PEATONAL_FILS <= NOT("0000000000010000");
					WHEN 6	 => PEATONAL_FILS <= NOT("0000000000100000");
					WHEN 7	 => PEATONAL_FILS <= NOT("0000000001000000");
					WHEN 8	 => PEATONAL_FILS <= NOT("0000000010000000");
					WHEN 9	 => PEATONAL_FILS <= NOT("0000000100000000");
					WHEN 10	 => PEATONAL_FILS <= NOT("0000001000000000");
					WHEN 11	 => PEATONAL_FILS <= NOT("0000010000000000");
					WHEN 12	 => PEATONAL_FILS <= NOT("0000100000000000");
					WHEN 13	 => PEATONAL_FILS <= NOT("0001000000000000");
					WHEN 14	 => PEATONAL_FILS <= NOT("0010000000000000");
					WHEN 15	 => PEATONAL_FILS <= NOT("0100000000000000");
					WHEN 16	 => PEATONAL_FILS <= NOT("1000000000000000");
					WHEN OTHERS	 => PEATONAL_FILS <= NOT("0000000000000000");
				END CASE;
				IF FILAS = 16 THEN FILAS <= 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	--PEATONAL--------------------------------------------
	PROCESS(CLK, CONTADOR, PEATONAL_FILS, ANIMACION) BEGIN
		IF RISING_EDGE(CLK) THEN
			IF ANIMACION = "00" THEN
				CASE PEATONAL_FILS IS
					WHEN "0000000000000001" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000000010" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000000100" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000001000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000010000" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000100000" 	=> PEATONAL_COLS <= "01111100";
					WHEN "0000000001000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000000010000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000000100000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000001000000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000010000000000" 	=> PEATONAL_COLS <= "10111000";
					WHEN "0000100000000000" 	=> PEATONAL_COLS <= "00111000";
					WHEN "0001000000000000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0010000000000000"		=> PEATONAL_COLS <= "00101000";
					WHEN "0100000000000000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "1000000000000000" 	=> PEATONAL_COLS <= "01111000";
					WHEN OTHERS => PEATONAL_COLS <= "00000000";
				END CASE;
			ELSIF ANIMACION = "01" THEN
				CASE PEATONAL_FILS IS
					WHEN "0000000000000001" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000000010" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000000100" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000001000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000010000" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000100000"		=> PEATONAL_COLS <= "01111100";
					WHEN "0000000001000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000000010000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000000100000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000001000000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000010000000000" 	=> PEATONAL_COLS <= "10111000";
					WHEN "0000100000000000" 	=> PEATONAL_COLS <= "00111000";
					WHEN "0001000000000000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0010000000000000" 	=> PEATONAL_COLS <= "00101110";
					WHEN "0100000000000000" 	=> PEATONAL_COLS <= "00100010";
					WHEN "1000000000000000" 	=> PEATONAL_COLS <= "01100000";
					WHEN OTHERS => PEATONAL_COLS <= "00000000";
				END CASE;
			ELSIF ANIMACION = "10" THEN
				CASE PEATONAL_FILS IS
					WHEN "0000000000000001"		=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000000010" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000000100" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000001000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000010000" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000100000" 	=> PEATONAL_COLS <= "01111100";
					WHEN "0000000001000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000000010000000" 	=> PEATONAL_COLS <= "01111001";
					WHEN "0000000100000000" 	=> PEATONAL_COLS <= "01111001";
					WHEN "0000001000000000" 	=> PEATONAL_COLS <= "11111001";
					WHEN "0000010000000000" 	=> PEATONAL_COLS <= "00111000";
					WHEN "0000100000000000" 	=> PEATONAL_COLS <= "00111000";
					WHEN "0001000000000000" 	=> PEATONAL_COLS <= "01001111";
					WHEN "0010000000000000" 	=> PEATONAL_COLS <= "01000001";
					WHEN "0100000000000000" 	=> PEATONAL_COLS <= "01000000";
					WHEN "1000000000000000" 	=> PEATONAL_COLS <= "11000000";
					WHEN OTHERS => PEATONAL_COLS <= "00000000";
				END CASE;
			ELSIF ANIMACION = "11" THEN
				CASE PEATONAL_FILS IS
					WHEN "0000000000000001" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000000010" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000000100" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000001000" 	=> PEATONAL_COLS <= "00101000";
					WHEN "0000000000010000" 	=> PEATONAL_COLS <= "00010000";
					WHEN "0000000000100000" 	=> PEATONAL_COLS <= "01111100";
					WHEN "0000000001000000" 	=> PEATONAL_COLS <= "01111010";
					WHEN "0000000010000000" 	=> PEATONAL_COLS <= "01111001";
					WHEN "0000000100000000" 	=> PEATONAL_COLS <= "01111001";
					WHEN "0000001000000000" 	=> PEATONAL_COLS <= "01111001";
					WHEN "0000010000000000" 	=> PEATONAL_COLS <= "10111000";
					WHEN "0000100000000000" 	=> PEATONAL_COLS <= "00111000";
					WHEN "0001000000000000" 	=> PEATONAL_COLS <= "11101000";
					WHEN "0010000000000000" 	=> PEATONAL_COLS <= "00001000";
					WHEN "0100000000000000" 	=> PEATONAL_COLS <= "00001000";
					WHEN "1000000000000000" 	=> PEATONAL_COLS <= "00011000";
					WHEN OTHERS => PEATONAL_COLS <= "00000000";
				END CASE;
			END IF;
		END IF;
	END PROCESS;
	
end Behavioral;

