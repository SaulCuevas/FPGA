`timescale 1ns / 1ps
//	INSTITUTO POLITECNICO NACIONAL
//					UPIITA
// AUTORES: SAUL CUEVAS MORALES
//				ALEXIS GONZALEZ ZUNIGA
// COMPARADOR DE MAGNITUD DE 4 BITS CON CODIFICADOR A DISPLAY Y BOTONES DE SELECTOR DE MODO
module P1_4bitMagnitudeComparator(
	
    );


endmodule
