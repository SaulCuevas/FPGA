----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SEMAFOROS is
end SEMAFOROS;

architecture Behavioral of SEMAFOROS is

begin


end Behavioral;

